`timescale 1ns / 1ps

module memory(//input
				clk,MemRead,MemWrite,IorD,IRWrite,
				PC,ALUOut,wdata,
				//output
				dataout,IR
    );
	input clk,MemRead,MemWrite,IorD,IRWrite;
	input[31:0] PC,ALUOut,wdata; //wdataΪ����д���ڴ������
	output[31:0] dataout;
	output reg[31:0] IR;
	
	wire[31:0] addr;

	assign addr=(IorD==0)?PC:ALUOut; //ѡ���ڴ���ʵ�ַ
	initial begin
		IR=0;
	end
	ram ram(
			.clka(clk),
			.addra(addr[8:0]),
			.dina(wdata),
			.douta(dataout),
			.wea(MemWrite)
			);

	always@*
	begin
		if(IRWrite==1)
			IR<=dataout; //дIR�Ĵ���
	end
endmodule
